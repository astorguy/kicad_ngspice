.title KiCad schematic
.tran 1n 300n
V2 vdc GND DC 2.345
R4 vpulse GND 10k
V5 vpwl GND pwl(0 -7 50n -7 51n -3 97n -4 171n -6.5 200n -6.5)
R1 vam GND 10k
R2 vdc GND 10k
R3 vexp GND 10k
V1 vam GND am(0.5 1 10meg 50meg 20n)
R6 vsffm GND 10k
R7 vsin GND 10k
R8 vtrnoise GND 10k
V6 vsffm GND sffm(-5 1 100meg 5 10meg)
V7 vsin GND DC 0 SIN( 0 1 100Meg 1n 10G )
R13 ipulse GND 10k
R14 ipwl GND 10k
I6 isffm GND sffm(-5 1 100meg 5 10meg)
I5 ipwl GND pwl(0 -7 50n -7 51n -3 97n -4 171n -6.5 200n -6.5)
R15 isffm GND 10k
I7 isin GND DC 0 SIN( 0 1 100Meg 1n 10G )
I1 iam GND am(0.5 1 10meg 50meg 20n)
I4 ipulse GND PULSE( -1 1 2n 30n 2n 50n 100n )
I3 iexp GND EXP( -4 -1 2n 30n 60n 40n )
R12 iexp GND 10k
R11 idc GND 10k
I2 idc GND DC 2.345
R10 iam GND 10k
V4 vpulse GND PULSE( -1 1 2n 30n 2n 50n 100n )
V3 vexp GND EXP( -4 -1 2n 30n 60n 40n )
R5 vpwl GND 10k
V9 vtrrandom GND TRRANDOM( 1 0 1 2 100n 98.000000 51.000000 )
R9 vtrrandom GND 10k
V8 vtrnoise GND TRNOISE( 100m 500p 0 0 0 0 0 ) AC 0 0
R18 itrrandom GND 10k
I9 itrrandom GND TRRANDOM( 1 0 1 2 100n 98.000000 51.000000 )
I8 itrnoise GND TRNOISE( 100m 500p 0 0 0 0 0 ) AC 0 0
R16 isin GND 10k
R17 itrnoise GND 10k
.end
