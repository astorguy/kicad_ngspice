.title KiCad schematic
.tran 10p 150n
V1 in GND PULSE( 0 3 100n 1n 1n 20n 100n )
R1 Net-_U1--_ GND 220
R2 Net-_U1-+_ in 160
C1 Net-_U1--_ Net-_Q1-E_ 1p
R3 Net-_Q1-E_ Net-_U1--_ 220
U1 Net-_U1-+_ Net-_U1--_ VDD VSS Net-_Q1-B_ __U1
Q1 VDD Net-_Q1-B_ Net-_Q1-E_ __Q1
R4 out Net-_U1-+_ 220
R5 out Net-_Q1-E_ 2.5
D1 out GND __D1
C2 out Net-_Q1-E_ 1p
V2 VDD GND DC 10
V3 GND VSS DC 10
.end
