.title KiCad schematic
.model Q2N2222 npn (bf=200)
.ac dec 100 10 1Meg

C4 VOUT Net-_C4-Pad2_ 10n
L1 Net-_C4-Pad2_ VOUT 100m
R1 +12V Net-_C4-Pad2_ 10
R2 VOUT Net-_C4-Pad2_ 22k
Q2 Net-_Q2-C_ VIN Net-_Q2-E_ Q2N2222
C2 VBASE 0 220p
Q1 VOUT VBASE Net-_Q1-E_ Q2N2222
R11 Net-_Q3-B_ 0 10k
R5 +12V VBASE 1k
R6 +12V Net-_Q3-B_ 22k
R3 +12V VIN 22k
R4 +12V Net-_Q2-C_ 1k
Q3 VBASE Net-_Q3-B_ Net-_Q2-E_ Q2N2222
R9 VIN 0 10k
R10 Net-_Q2-E_ 0 470
C1 VIN Net-_V2-E1_ 1U
V2 Net-_V2-E1_ 0 dc 0 ac 1
V1 +12V 0 DC 12
R8 Net-_Q1-E_ 0 2.2k
R12 Net-_L2-Pad1_ Net-_Q1-E_ 100
R7 Net-_C3-Pad1_ Net-_L2-Pad1_ 22k
L2 Net-_L2-Pad1_ Net-_C3-Pad1_ 100m
C3 Net-_C3-Pad1_ 0 10n
.end
