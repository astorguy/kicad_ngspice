.title KiCad schematic
.include "/workspaces/kicad_ngspice/examples/from_kicad_distribution/sallen_key/ad8051.lib"
.control
version
.endc
.ac dec 10 1 1Meg

C2 Net-_U1-+_ GND 100n
R2 Net-_U1-+_ Net-_C1-Pad2_ 1k
R1 Net-_C1-Pad2_ Net-_R1-Pad2_ 1k
V1 Net-_R1-Pad2_ GND ac=1
C1 lowpass Net-_C1-Pad2_ 100n
XU1 Net-_U1-+_ lowpass VDD VSS lowpass AD8051
V2 VDD GND DC 10
V3 GND VSS DC 10
.end
